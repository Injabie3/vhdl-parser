Library ieee;Use ieee.std_logic_1164.all;Use ieee.numeric_std.all;Entity Over60 isPORT (    X     : IN unsigned(5 DOWNTO 0);    Y    : OUT std_logic);End Entity Over60;Architecture behavior of Over60 isBeginY <= (X(5) AND X(4) AND X(3) AND X(2)) after 8 ns; -- COMMENT When the four leftmost bits are 1 then the number is over 60End Architecture behavior;--The comment at the end.