'0' '1'
'-' 'z'
